///////////////////////////////////////////////////////////////////////////////////////////////////
//
// UVM SPI MEM TB pkg
// 
// This is the top level SPIMEM testbench package 
// SPI MEM
//
///////////////////////////////////////////////////////////////////////////////////////////////////

 package SPI_Mem_TB_pkg;
 
  import UVM_SPI_Mem_TB_Tests_pkg::*;
  
 endpackage