
//==============================================================
// File: UVM_SPI_Mem_TB_pkg.sv
// Description: SPI Agent Package - SPI-MEMORY.
//
// Author: Grupo de Verificación
//==============================================================

